module dataMemory (address,write_data, memwrite, memread,clk,read_data );
parameter Width = 32;
input  [Width-1:0] address; 
input  [Width-1:0] write_data;    
input  memwrite, memread,clk;         
output reg [Width-1:0] read_data;   
reg [Width-1:0] mem [0:255]; 

integer i;

initial begin
  read_data <= 0;
  for (i = 0; i < 256; i = i + 1) begin
    mem[i] = i;
  end
end

always @(posedge clk) begin
  if (memwrite == 1'b1) begin
    mem[address] <= write_data;
  end
 
  if (memread == 1'b1) begin
    read_data <= mem[address];
  end
end

endmodule