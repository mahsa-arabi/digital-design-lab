module clock (clk);
output reg clk;
                    
initial begin
        clk = 1'b0;
end
endmodule